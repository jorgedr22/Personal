timescale 1ns/1ps

module EX3 (go,done,min,sum,CLK,Rst);
    input go, CLK, Rst;
    output reg done;
    output reg [8:0] min, sum;

    







endmodule